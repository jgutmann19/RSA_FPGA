// // This module computes m^e % n
module modexp #(
    parameter int WIDTH
)(
    input
);

endmodule